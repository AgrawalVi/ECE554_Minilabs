// Deprecated file kept for compatibility with prior lab checkouts.
// Use matrix_vector_multi.sv (underscore) instead.
